module top #(
  parameter int XLEN = 32
) (
  input logic clk,
  input logic n_rst
);

endmodule
