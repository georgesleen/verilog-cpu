parameter int XLEN = 32;
